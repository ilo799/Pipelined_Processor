module Testbench;
endmodule
//Testbenches don't have ports

