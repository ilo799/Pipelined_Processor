module Processor (clk, reset);
 input clk, reset;
endmodule
